`ifndef RAM_V_ 
`define RAM_V_ 

module RAM(
    
);
endmodule

`endif